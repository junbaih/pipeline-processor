`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 01/07/2018 10:21:50 PM
// Design Name: 
// Module Name: mux2
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mux2
    #(parameter WIDTH = 32)
    (input logic [WIDTH-1:0] d0, d1,d2,d3,d4,
     input logic [2:0] s,
     output logic [WIDTH-1:0] y);

assign y = s==3'b0 ? d0 : (s==3'b001?d1:(s==3'b010?d2:(s==3'b011?d3:d4)));

endmodule
